/*
Assignment: A21

Update code mentioned in the Instruction tab to send your name on Console. 
*/

`include "uvm_macros.svh"
import uvm_pkg::*;  //compiler directives

module tb;
  
  initial begin
    `uvm_info("TB_TOP", "SAIKRUPA", UVM_MEDIUM); //id, msg, verbosity level
  end
  
endmodule